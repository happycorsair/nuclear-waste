/* Definition of the `ping` component. */

component mosquitto.Ping

endpoints {
    /* Declaration of a named implementation of the "Ping" interface. */
    ping : mosquitto.Ping
}
